// 0716089
//Subject:      CO project 2 - Shift_Left_Two_32
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Description: 
//--------------------------------------------------------------------------------
`timescale 1ns/1ps
module Shift_Left_Two_32(
    data_i,
    data_o
    );

//I/O ports                    
input [32-1:0] data_i;
output [32-1:0] data_o;
reg[32-1:0] data_o;
wire[32-1:0] temp;
assign temp = data_i << 2;
//shift left 2
always @(*) begin
    data_o = temp;
end
endmodule
